module MY_BUS(
		
		);

endmodule
