`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:45:58 07/21/2016 
// Design Name: 
// Module Name:    charvram_mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module charvram_mux(
	input reg [12:0] addr_cpu,
	input reg [7:0] data_cpu,
	input reg wea,
	
	input
    );

endmodule
